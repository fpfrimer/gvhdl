---------------------------------------------------
-- File: <entity_name>.vhd
-- Developer: developer_name
-- Company: company_name
-- Date: <date>
---------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity <entity_name> is
    port (
        -- list of input/output ports
        <port_list>
    );
end <entity_name>;

architecture <architecture_name> of <entity_name> is
    -- signal, component declarations, etc.
begin
    -- circuit behavior description
end <architecture_name>;